// Copyright 2021 
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
// Licensed under the Solderpad Hardware License v 2.1 (the "License"); you may not use this file except in compliance
// with the License, or, at your option, the Apache License version 2.0.  You may obtain a copy of the License at
//                                        https://solderpad.org/licenses/SHL-2.1/
// Unless required by applicable law or agreed to in writing, any work distributed under the License is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.  See the License for the
// specific language governing permissions and limitations under the License.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_DP_CHKR_SV__
`define __UVME_DP_CHKR_SV__


/**
 * TODO Describe uvme_dp_chkr
 */
module uvme_dp_chkr (
   // TODO Add interfaces to uvme_dp_chkr
);
   
   // TODO Add assertions to uvme_$[name}_chkr
   
endmodule : uvme_dp_chkr


`endif // __UVME_DP_CHKR_SV__
